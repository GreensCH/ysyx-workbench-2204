`timescale 1ps/1ps
module rom_ps2kbd_ascii(
	input   [7:0]     addr,
	output reg [7:0]    data
);
    always@(*)begin
        case(addr)
            8'h0E:data=8'h60;//~
            8'h16:data=8'h31;//1
            8'h1E:data=8'h32;//2
            8'h26:data=8'h33;//3
            8'h25:data=8'h34;//4
            8'h2E:data=8'h35;//5
            8'h36:data=8'h36;//6
            8'h3D:data=8'h37;//7
            8'h3E:data=8'h38;//8
            8'h46:data=8'h39;//9
            8'h45:data=8'h30;//0
            8'h4E:data=8'h2D;//-
            8'h55:data=8'h3D;//=
            8'h1C:data=8'h61;//a
            8'h32:data=8'h62;//b
            8'h21:data=8'h63;//c
            8'h23:data=8'h64;//d
            8'h24:data=8'h65;//e
            8'h2B:data=8'h66;//f
            8'h34:data=8'h67;//g
            8'h33:data=8'h68;//h
            8'h43:data=8'h69;//i
            8'h3B:data=8'h6A;//j
            8'h42:data=8'h6B;//k
            8'h4B:data=8'h6C;//l
            8'h3A:data=8'h6D;//m
            8'h31:data=8'h6E;//n
            8'h44:data=8'h6F;//o
            8'h4D:data=8'h70;//p
            8'h15:data=8'h71;//q
            8'h2D:data=8'h72;//r
            8'h1B:data=8'h73;//s
            8'h2C:data=8'h74;//t
            8'h3C:data=8'h75;//u
            8'h2A:data=8'h76;//v
            8'h1D:data=8'h77;//w
            8'h22:data=8'h78;//x
            8'h35:data=8'h79;//y
            8'h1A:data=8'h7A;//z
            8'h0D:data=8'd09;//TAB
            8'h58:data=8'd20;//Caps?
            8'h12:data=8'd16;//Shift?
            8'h14:data=8'd17;//Ctrl?
            8'h11:data=8'd18;//Alt?
            8'h29:data=8'd32;//space
            8'h54:data=8'd219;//[
            8'h5B:data=8'd221;//]
            8'h5D:data=8'd220;//\|
            8'h4C:data=8'd186;//;
            8'h52:data=8'd222;//“
            8'h41:data=8'd220;//，<
            8'h49:data=8'd110;//.>
            8'h6B:data=8'd37;//left
            8'h75:data=8'd38;//up
            8'h74:data=8'd39;//right
            8'h72:data=8'd40;//down
            8'h71:data=8'd46;//delete
            8'h77:data=8'd144;//num lock
            8'h66:data=8'd08;//backspcase
            8'h76:data=8'd27;//escape
            8'h05:data=8'd112;//F1
            8'h06:data=8'd113;//F2
            8'h04:data=8'd114;//F3
            8'h0C:data=8'd115;//F4
            8'h03:data=8'd116;//F5
            8'h0B:data=8'd117;//F6
            8'h83:data=8'd118;//F7
            8'h0A:data=8'd119;//F8
            8'h01:data=8'd120;//F8
            8'h09:data=8'd121;//F9
            8'h78:data=8'd122;//F10
            8'h07:data=8'd123;//F11
            default:data=8'h0;
        endcase
    end

endmodule